module mult(
    input  wire        mul_clk    ,
    input  wire        rst        ,
    input  wire        mul        ,
    input  wire        mul_signed ,
    input  wire [31:0] x          ,
    input  wire [31:0] y          ,
    output reg  [63:0] result     ,
    output wire        complete
);

integer i;
assign complete = i;
always @(posedge mul_clk) begin
        i<= rst ? 0: (i == 1)? 0: (mul) ? i + 1 : i;
end

always @(posedge mul_clk) begin
    if(rst)
        result <= 0;
    else
        result <= P[63:0];    
end


wire [32:0] A = ({{ mul_signed & x[31]}, x})
              | ({{!mul_signed & 1'b0 }, x});
wire [32:0] B = ({{ mul_signed & y[31]}, y})
              | ({{!mul_signed & 1'b0 }, y});

wire [65:0] p00, p01, p02, p03, p04, p05, p06, p07, p08, p09, p10, p11, p12, p13, p14, p15, p16;
wire        C00, C01, C02, C03, C04, C05, C06, C07, C08, C09, C10, C11, C12, C13, C14, C15, C16;

wire [65:0] S, C;

wire [65:0] P = S + {C[64:0], C15} + {65'd0, C16};

wire [16:0] s00 = {p16[ 0], p15[ 0], p14[ 0], p13[ 0], p12[ 0], p11[ 0], p10[ 0], p09[ 0], p08[ 0], p07[ 0], p06[ 0], p05[ 0], p04[ 0], p03[ 0], p02[ 0], p01[ 0], p00[ 0]};
wire [16:0] s01 = {p16[ 1], p15[ 1], p14[ 1], p13[ 1], p12[ 1], p11[ 1], p10[ 1], p09[ 1], p08[ 1], p07[ 1], p06[ 1], p05[ 1], p04[ 1], p03[ 1], p02[ 1], p01[ 1], p00[ 1]};
wire [16:0] s02 = {p16[ 2], p15[ 2], p14[ 2], p13[ 2], p12[ 2], p11[ 2], p10[ 2], p09[ 2], p08[ 2], p07[ 2], p06[ 2], p05[ 2], p04[ 2], p03[ 2], p02[ 2], p01[ 2], p00[ 2]};
wire [16:0] s03 = {p16[ 3], p15[ 3], p14[ 3], p13[ 3], p12[ 3], p11[ 3], p10[ 3], p09[ 3], p08[ 3], p07[ 3], p06[ 3], p05[ 3], p04[ 3], p03[ 3], p02[ 3], p01[ 3], p00[ 3]};
wire [16:0] s04 = {p16[ 4], p15[ 4], p14[ 4], p13[ 4], p12[ 4], p11[ 4], p10[ 4], p09[ 4], p08[ 4], p07[ 4], p06[ 4], p05[ 4], p04[ 4], p03[ 4], p02[ 4], p01[ 4], p00[ 4]};
wire [16:0] s05 = {p16[ 5], p15[ 5], p14[ 5], p13[ 5], p12[ 5], p11[ 5], p10[ 5], p09[ 5], p08[ 5], p07[ 5], p06[ 5], p05[ 5], p04[ 5], p03[ 5], p02[ 5], p01[ 5], p00[ 5]};
wire [16:0] s06 = {p16[ 6], p15[ 6], p14[ 6], p13[ 6], p12[ 6], p11[ 6], p10[ 6], p09[ 6], p08[ 6], p07[ 6], p06[ 6], p05[ 6], p04[ 6], p03[ 6], p02[ 6], p01[ 6], p00[ 6]};
wire [16:0] s07 = {p16[ 7], p15[ 7], p14[ 7], p13[ 7], p12[ 7], p11[ 7], p10[ 7], p09[ 7], p08[ 7], p07[ 7], p06[ 7], p05[ 7], p04[ 7], p03[ 7], p02[ 7], p01[ 7], p00[ 7]};
wire [16:0] s08 = {p16[ 8], p15[ 8], p14[ 8], p13[ 8], p12[ 8], p11[ 8], p10[ 8], p09[ 8], p08[ 8], p07[ 8], p06[ 8], p05[ 8], p04[ 8], p03[ 8], p02[ 8], p01[ 8], p00[ 8]};
wire [16:0] s09 = {p16[ 9], p15[ 9], p14[ 9], p13[ 9], p12[ 9], p11[ 9], p10[ 9], p09[ 9], p08[ 9], p07[ 9], p06[ 9], p05[ 9], p04[ 9], p03[ 9], p02[ 9], p01[ 9], p00[ 9]};
wire [16:0] s10 = {p16[10], p15[10], p14[10], p13[10], p12[10], p11[10], p10[10], p09[10], p08[10], p07[10], p06[10], p05[10], p04[10], p03[10], p02[10], p01[10], p00[10]};
wire [16:0] s11 = {p16[11], p15[11], p14[11], p13[11], p12[11], p11[11], p10[11], p09[11], p08[11], p07[11], p06[11], p05[11], p04[11], p03[11], p02[11], p01[11], p00[11]};
wire [16:0] s12 = {p16[12], p15[12], p14[12], p13[12], p12[12], p11[12], p10[12], p09[12], p08[12], p07[12], p06[12], p05[12], p04[12], p03[12], p02[12], p01[12], p00[12]};
wire [16:0] s13 = {p16[13], p15[13], p14[13], p13[13], p12[13], p11[13], p10[13], p09[13], p08[13], p07[13], p06[13], p05[13], p04[13], p03[13], p02[13], p01[13], p00[13]};
wire [16:0] s14 = {p16[14], p15[14], p14[14], p13[14], p12[14], p11[14], p10[14], p09[14], p08[14], p07[14], p06[14], p05[14], p04[14], p03[14], p02[14], p01[14], p00[14]};
wire [16:0] s15 = {p16[15], p15[15], p14[15], p13[15], p12[15], p11[15], p10[15], p09[15], p08[15], p07[15], p06[15], p05[15], p04[15], p03[15], p02[15], p01[15], p00[15]};
wire [16:0] s16 = {p16[16], p15[16], p14[16], p13[16], p12[16], p11[16], p10[16], p09[16], p08[16], p07[16], p06[16], p05[16], p04[16], p03[16], p02[16], p01[16], p00[16]};
wire [16:0] s17 = {p16[17], p15[17], p14[17], p13[17], p12[17], p11[17], p10[17], p09[17], p08[17], p07[17], p06[17], p05[17], p04[17], p03[17], p02[17], p01[17], p00[17]};
wire [16:0] s18 = {p16[18], p15[18], p14[18], p13[18], p12[18], p11[18], p10[18], p09[18], p08[18], p07[18], p06[18], p05[18], p04[18], p03[18], p02[18], p01[18], p00[18]};
wire [16:0] s19 = {p16[19], p15[19], p14[19], p13[19], p12[19], p11[19], p10[19], p09[19], p08[19], p07[19], p06[19], p05[19], p04[19], p03[19], p02[19], p01[19], p00[19]};
wire [16:0] s20 = {p16[20], p15[20], p14[20], p13[20], p12[20], p11[20], p10[20], p09[20], p08[20], p07[20], p06[20], p05[20], p04[20], p03[20], p02[20], p01[20], p00[20]};
wire [16:0] s21 = {p16[21], p15[21], p14[21], p13[21], p12[21], p11[21], p10[21], p09[21], p08[21], p07[21], p06[21], p05[21], p04[21], p03[21], p02[21], p01[21], p00[21]};
wire [16:0] s22 = {p16[22], p15[22], p14[22], p13[22], p12[22], p11[22], p10[22], p09[22], p08[22], p07[22], p06[22], p05[22], p04[22], p03[22], p02[22], p01[22], p00[22]};
wire [16:0] s23 = {p16[23], p15[23], p14[23], p13[23], p12[23], p11[23], p10[23], p09[23], p08[23], p07[23], p06[23], p05[23], p04[23], p03[23], p02[23], p01[23], p00[23]};
wire [16:0] s24 = {p16[24], p15[24], p14[24], p13[24], p12[24], p11[24], p10[24], p09[24], p08[24], p07[24], p06[24], p05[24], p04[24], p03[24], p02[24], p01[24], p00[24]};
wire [16:0] s25 = {p16[25], p15[25], p14[25], p13[25], p12[25], p11[25], p10[25], p09[25], p08[25], p07[25], p06[25], p05[25], p04[25], p03[25], p02[25], p01[25], p00[25]};
wire [16:0] s26 = {p16[26], p15[26], p14[26], p13[26], p12[26], p11[26], p10[26], p09[26], p08[26], p07[26], p06[26], p05[26], p04[26], p03[26], p02[26], p01[26], p00[26]};
wire [16:0] s27 = {p16[27], p15[27], p14[27], p13[27], p12[27], p11[27], p10[27], p09[27], p08[27], p07[27], p06[27], p05[27], p04[27], p03[27], p02[27], p01[27], p00[27]};
wire [16:0] s28 = {p16[28], p15[28], p14[28], p13[28], p12[28], p11[28], p10[28], p09[28], p08[28], p07[28], p06[28], p05[28], p04[28], p03[28], p02[28], p01[28], p00[28]};
wire [16:0] s29 = {p16[29], p15[29], p14[29], p13[29], p12[29], p11[29], p10[29], p09[29], p08[29], p07[29], p06[29], p05[29], p04[29], p03[29], p02[29], p01[29], p00[29]};
wire [16:0] s30 = {p16[30], p15[30], p14[30], p13[30], p12[30], p11[30], p10[30], p09[30], p08[30], p07[30], p06[30], p05[30], p04[30], p03[30], p02[30], p01[30], p00[30]};
wire [16:0] s31 = {p16[31], p15[31], p14[31], p13[31], p12[31], p11[31], p10[31], p09[31], p08[31], p07[31], p06[31], p05[31], p04[31], p03[31], p02[31], p01[31], p00[31]};
wire [16:0] s32 = {p16[32], p15[32], p14[32], p13[32], p12[32], p11[32], p10[32], p09[32], p08[32], p07[32], p06[32], p05[32], p04[32], p03[32], p02[32], p01[32], p00[32]};
wire [16:0] s33 = {p16[33], p15[33], p14[33], p13[33], p12[33], p11[33], p10[33], p09[33], p08[33], p07[33], p06[33], p05[33], p04[33], p03[33], p02[33], p01[33], p00[33]};
wire [16:0] s34 = {p16[34], p15[34], p14[34], p13[34], p12[34], p11[34], p10[34], p09[34], p08[34], p07[34], p06[34], p05[34], p04[34], p03[34], p02[34], p01[34], p00[34]};
wire [16:0] s35 = {p16[35], p15[35], p14[35], p13[35], p12[35], p11[35], p10[35], p09[35], p08[35], p07[35], p06[35], p05[35], p04[35], p03[35], p02[35], p01[35], p00[35]};
wire [16:0] s36 = {p16[36], p15[36], p14[36], p13[36], p12[36], p11[36], p10[36], p09[36], p08[36], p07[36], p06[36], p05[36], p04[36], p03[36], p02[36], p01[36], p00[36]};
wire [16:0] s37 = {p16[37], p15[37], p14[37], p13[37], p12[37], p11[37], p10[37], p09[37], p08[37], p07[37], p06[37], p05[37], p04[37], p03[37], p02[37], p01[37], p00[37]};
wire [16:0] s38 = {p16[38], p15[38], p14[38], p13[38], p12[38], p11[38], p10[38], p09[38], p08[38], p07[38], p06[38], p05[38], p04[38], p03[38], p02[38], p01[38], p00[38]};
wire [16:0] s39 = {p16[39], p15[39], p14[39], p13[39], p12[39], p11[39], p10[39], p09[39], p08[39], p07[39], p06[39], p05[39], p04[39], p03[39], p02[39], p01[39], p00[39]};
wire [16:0] s40 = {p16[40], p15[40], p14[40], p13[40], p12[40], p11[40], p10[40], p09[40], p08[40], p07[40], p06[40], p05[40], p04[40], p03[40], p02[40], p01[40], p00[40]};
wire [16:0] s41 = {p16[41], p15[41], p14[41], p13[41], p12[41], p11[41], p10[41], p09[41], p08[41], p07[41], p06[41], p05[41], p04[41], p03[41], p02[41], p01[41], p00[41]};
wire [16:0] s42 = {p16[42], p15[42], p14[42], p13[42], p12[42], p11[42], p10[42], p09[42], p08[42], p07[42], p06[42], p05[42], p04[42], p03[42], p02[42], p01[42], p00[42]};
wire [16:0] s43 = {p16[43], p15[43], p14[43], p13[43], p12[43], p11[43], p10[43], p09[43], p08[43], p07[43], p06[43], p05[43], p04[43], p03[43], p02[43], p01[43], p00[43]};
wire [16:0] s44 = {p16[44], p15[44], p14[44], p13[44], p12[44], p11[44], p10[44], p09[44], p08[44], p07[44], p06[44], p05[44], p04[44], p03[44], p02[44], p01[44], p00[44]};
wire [16:0] s45 = {p16[45], p15[45], p14[45], p13[45], p12[45], p11[45], p10[45], p09[45], p08[45], p07[45], p06[45], p05[45], p04[45], p03[45], p02[45], p01[45], p00[45]};
wire [16:0] s46 = {p16[46], p15[46], p14[46], p13[46], p12[46], p11[46], p10[46], p09[46], p08[46], p07[46], p06[46], p05[46], p04[46], p03[46], p02[46], p01[46], p00[46]};
wire [16:0] s47 = {p16[47], p15[47], p14[47], p13[47], p12[47], p11[47], p10[47], p09[47], p08[47], p07[47], p06[47], p05[47], p04[47], p03[47], p02[47], p01[47], p00[47]};
wire [16:0] s48 = {p16[48], p15[48], p14[48], p13[48], p12[48], p11[48], p10[48], p09[48], p08[48], p07[48], p06[48], p05[48], p04[48], p03[48], p02[48], p01[48], p00[48]};
wire [16:0] s49 = {p16[49], p15[49], p14[49], p13[49], p12[49], p11[49], p10[49], p09[49], p08[49], p07[49], p06[49], p05[49], p04[49], p03[49], p02[49], p01[49], p00[49]};
wire [16:0] s50 = {p16[50], p15[50], p14[50], p13[50], p12[50], p11[50], p10[50], p09[50], p08[50], p07[50], p06[50], p05[50], p04[50], p03[50], p02[50], p01[50], p00[50]};
wire [16:0] s51 = {p16[51], p15[51], p14[51], p13[51], p12[51], p11[51], p10[51], p09[51], p08[51], p07[51], p06[51], p05[51], p04[51], p03[51], p02[51], p01[51], p00[51]};
wire [16:0] s52 = {p16[52], p15[52], p14[52], p13[52], p12[52], p11[52], p10[52], p09[52], p08[52], p07[52], p06[52], p05[52], p04[52], p03[52], p02[52], p01[52], p00[52]};
wire [16:0] s53 = {p16[53], p15[53], p14[53], p13[53], p12[53], p11[53], p10[53], p09[53], p08[53], p07[53], p06[53], p05[53], p04[53], p03[53], p02[53], p01[53], p00[53]};
wire [16:0] s54 = {p16[54], p15[54], p14[54], p13[54], p12[54], p11[54], p10[54], p09[54], p08[54], p07[54], p06[54], p05[54], p04[54], p03[54], p02[54], p01[54], p00[54]};
wire [16:0] s55 = {p16[55], p15[55], p14[55], p13[55], p12[55], p11[55], p10[55], p09[55], p08[55], p07[55], p06[55], p05[55], p04[55], p03[55], p02[55], p01[55], p00[55]};
wire [16:0] s56 = {p16[56], p15[56], p14[56], p13[56], p12[56], p11[56], p10[56], p09[56], p08[56], p07[56], p06[56], p05[56], p04[56], p03[56], p02[56], p01[56], p00[56]};
wire [16:0] s57 = {p16[57], p15[57], p14[57], p13[57], p12[57], p11[57], p10[57], p09[57], p08[57], p07[57], p06[57], p05[57], p04[57], p03[57], p02[57], p01[57], p00[57]};
wire [16:0] s58 = {p16[58], p15[58], p14[58], p13[58], p12[58], p11[58], p10[58], p09[58], p08[58], p07[58], p06[58], p05[58], p04[58], p03[58], p02[58], p01[58], p00[58]};
wire [16:0] s59 = {p16[59], p15[59], p14[59], p13[59], p12[59], p11[59], p10[59], p09[59], p08[59], p07[59], p06[59], p05[59], p04[59], p03[59], p02[59], p01[59], p00[59]};
wire [16:0] s60 = {p16[60], p15[60], p14[60], p13[60], p12[60], p11[60], p10[60], p09[60], p08[60], p07[60], p06[60], p05[60], p04[60], p03[60], p02[60], p01[60], p00[60]};
wire [16:0] s61 = {p16[61], p15[61], p14[61], p13[61], p12[61], p11[61], p10[61], p09[61], p08[61], p07[61], p06[61], p05[61], p04[61], p03[61], p02[61], p01[61], p00[61]};
wire [16:0] s62 = {p16[62], p15[62], p14[62], p13[62], p12[62], p11[62], p10[62], p09[62], p08[62], p07[62], p06[62], p05[62], p04[62], p03[62], p02[62], p01[62], p00[62]};
wire [16:0] s63 = {p16[63], p15[63], p14[63], p13[63], p12[63], p11[63], p10[63], p09[63], p08[63], p07[63], p06[63], p05[63], p04[63], p03[63], p02[63], p01[63], p00[63]};
wire [16:0] s64 = {p16[64], p15[64], p14[64], p13[64], p12[64], p11[64], p10[64], p09[64], p08[64], p07[64], p06[64], p05[64], p04[64], p03[64], p02[64], p01[64], p00[64]};
wire [16:0] s65 = {p16[65], p15[65], p14[65], p13[65], p12[65], p11[65], p10[65], p09[65], p08[65], p07[65], p06[65], p05[65], p04[65], p03[65], p02[65], p01[65], p00[65]};

wire [66:0] w00, w01, w02, w03, w04, w05, w06, w07, w08, w09, w10, w11, w12, w13, w14;

assign {w00[0],w01[0],w02[0],w03[0],w04[0],w05[0],w06[0],w07[0],w08[0],w09[0],w10[0],w11[0],w12[0],w13[0],w14[0]} 
     = {C00   ,C01   ,C02   ,C03   ,C04   ,C05   ,C06   ,C07   ,C08   ,C09   ,C10   ,C11   ,C12   ,C13   ,C14   };

mips_wallace_unit wallace_unit00(s00, w00[ 0], w01[ 0], w02[ 0], w03[ 0], w04[ 0], w05[ 0], w06[ 0], w07[ 0], w08[ 0], w09[ 0], w10[ 0], w11[ 0], w12[ 0], w13[ 0], w14[ 0],
                                      w00[ 1], w01[ 1], w02[ 1], w03[ 1], w04[ 1], w05[ 1], w06[ 1], w07[ 1], w08[ 1], w09[ 1], w10[ 1], w11[ 1], w12[ 1], w13[ 1], w14[ 1],
                                        S[ 0],   C[ 0]);
mips_wallace_unit wallace_unit01(s01, w00[ 1], w01[ 1], w02[ 1], w03[ 1], w04[ 1], w05[ 1], w06[ 1], w07[ 1], w08[ 1], w09[ 1], w10[ 1], w11[ 1], w12[ 1], w13[ 1], w14[ 1],
                                      w00[ 2], w01[ 2], w02[ 2], w03[ 2], w04[ 2], w05[ 2], w06[ 2], w07[ 2], w08[ 2], w09[ 2], w10[ 2], w11[ 2], w12[ 2], w13[ 2], w14[ 2],
                                        S[ 1],   C[ 1]);
mips_wallace_unit wallace_unit02(s02, w00[ 2], w01[ 2], w02[ 2], w03[ 2], w04[ 2], w05[ 2], w06[ 2], w07[ 2], w08[ 2], w09[ 2], w10[ 2], w11[ 2], w12[ 2], w13[ 2], w14[ 2],
                                      w00[ 3], w01[ 3], w02[ 3], w03[ 3], w04[ 3], w05[ 3], w06[ 3], w07[ 3], w08[ 3], w09[ 3], w10[ 3], w11[ 3], w12[ 3], w13[ 3], w14[ 3],
                                        S[ 2],   C[ 2]);
mips_wallace_unit wallace_unit03(s03, w00[ 3], w01[ 3], w02[ 3], w03[ 3], w04[ 3], w05[ 3], w06[ 3], w07[ 3], w08[ 3], w09[ 3], w10[ 3], w11[ 3], w12[ 3], w13[ 3], w14[ 3],
                                      w00[ 4], w01[ 4], w02[ 4], w03[ 4], w04[ 4], w05[ 4], w06[ 4], w07[ 4], w08[ 4], w09[ 4], w10[ 4], w11[ 4], w12[ 4], w13[ 4], w14[ 4],
                                        S[ 3],   C[ 3]);
mips_wallace_unit wallace_unit04(s04, w00[ 4], w01[ 4], w02[ 4], w03[ 4], w04[ 4], w05[ 4], w06[ 4], w07[ 4], w08[ 4], w09[ 4], w10[ 4], w11[ 4], w12[ 4], w13[ 4], w14[ 4],
                                      w00[ 5], w01[ 5], w02[ 5], w03[ 5], w04[ 5], w05[ 5], w06[ 5], w07[ 5], w08[ 5], w09[ 5], w10[ 5], w11[ 5], w12[ 5], w13[ 5], w14[ 5],
                                        S[ 4],   C[ 4]);
mips_wallace_unit wallace_unit05(s05, w00[ 5], w01[ 5], w02[ 5], w03[ 5], w04[ 5], w05[ 5], w06[ 5], w07[ 5], w08[ 5], w09[ 5], w10[ 5], w11[ 5], w12[ 5], w13[ 5], w14[ 5],
                                      w00[ 6], w01[ 6], w02[ 6], w03[ 6], w04[ 6], w05[ 6], w06[ 6], w07[ 6], w08[ 6], w09[ 6], w10[ 6], w11[ 6], w12[ 6], w13[ 6], w14[ 6],
                                        S[ 5],   C[ 5]);
mips_wallace_unit wallace_unit06(s06, w00[ 6], w01[ 6], w02[ 6], w03[ 6], w04[ 6], w05[ 6], w06[ 6], w07[ 6], w08[ 6], w09[ 6], w10[ 6], w11[ 6], w12[ 6], w13[ 6], w14[ 6],
                                      w00[ 7], w01[ 7], w02[ 7], w03[ 7], w04[ 7], w05[ 7], w06[ 7], w07[ 7], w08[ 7], w09[ 7], w10[ 7], w11[ 7], w12[ 7], w13[ 7], w14[ 7],
                                        S[ 6],   C[ 6]);
mips_wallace_unit wallace_unit07(s07, w00[ 7], w01[ 7], w02[ 7], w03[ 7], w04[ 7], w05[ 7], w06[ 7], w07[ 7], w08[ 7], w09[ 7], w10[ 7], w11[ 7], w12[ 7], w13[ 7], w14[ 7],
                                      w00[ 8], w01[ 8], w02[ 8], w03[ 8], w04[ 8], w05[ 8], w06[ 8], w07[ 8], w08[ 8], w09[ 8], w10[ 8], w11[ 8], w12[ 8], w13[ 8], w14[ 8],
                                        S[ 7],   C[ 7]);
mips_wallace_unit wallace_unit08(s08, w00[ 8], w01[ 8], w02[ 8], w03[ 8], w04[ 8], w05[ 8], w06[ 8], w07[ 8], w08[ 8], w09[ 8], w10[ 8], w11[ 8], w12[ 8], w13[ 8], w14[ 8],
                                      w00[ 9], w01[ 9], w02[ 9], w03[ 9], w04[ 9], w05[ 9], w06[ 9], w07[ 9], w08[ 9], w09[ 9], w10[ 9], w11[ 9], w12[ 9], w13[ 9], w14[ 9],
                                        S[ 8],   C[ 8]);
mips_wallace_unit wallace_unit09(s09, w00[ 9], w01[ 9], w02[ 9], w03[ 9], w04[ 9], w05[ 9], w06[ 9], w07[ 9], w08[ 9], w09[ 9], w10[ 9], w11[ 9], w12[ 9], w13[ 9], w14[ 9],
                                      w00[10], w01[10], w02[10], w03[10], w04[10], w05[10], w06[10], w07[10], w08[10], w09[10], w10[10], w11[10], w12[10], w13[10], w14[10],
                                        S[ 9],   C[ 9]);
mips_wallace_unit wallace_unit10(s10, w00[10], w01[10], w02[10], w03[10], w04[10], w05[10], w06[10], w07[10], w08[10], w09[10], w10[10], w11[10], w12[10], w13[10], w14[10],
                                      w00[11], w01[11], w02[11], w03[11], w04[11], w05[11], w06[11], w07[11], w08[11], w09[11], w10[11], w11[11], w12[11], w13[11], w14[11],
                                        S[10],   C[10]);
mips_wallace_unit wallace_unit11(s11, w00[11], w01[11], w02[11], w03[11], w04[11], w05[11], w06[11], w07[11], w08[11], w09[11], w10[11], w11[11], w12[11], w13[11], w14[11],
                                      w00[12], w01[12], w02[12], w03[12], w04[12], w05[12], w06[12], w07[12], w08[12], w09[12], w10[12], w11[12], w12[12], w13[12], w14[12],
                                        S[11],   C[11]);
mips_wallace_unit wallace_unit12(s12, w00[12], w01[12], w02[12], w03[12], w04[12], w05[12], w06[12], w07[12], w08[12], w09[12], w10[12], w11[12], w12[12], w13[12], w14[12],
                                      w00[13], w01[13], w02[13], w03[13], w04[13], w05[13], w06[13], w07[13], w08[13], w09[13], w10[13], w11[13], w12[13], w13[13], w14[13],
                                        S[12],   C[12]);
mips_wallace_unit wallace_unit13(s13, w00[13], w01[13], w02[13], w03[13], w04[13], w05[13], w06[13], w07[13], w08[13], w09[13], w10[13], w11[13], w12[13], w13[13], w14[13],
                                      w00[14], w01[14], w02[14], w03[14], w04[14], w05[14], w06[14], w07[14], w08[14], w09[14], w10[14], w11[14], w12[14], w13[14], w14[14],
                                        S[13],   C[13]);
mips_wallace_unit wallace_unit14(s14, w00[14], w01[14], w02[14], w03[14], w04[14], w05[14], w06[14], w07[14], w08[14], w09[14], w10[14], w11[14], w12[14], w13[14], w14[14],
                                      w00[15], w01[15], w02[15], w03[15], w04[15], w05[15], w06[15], w07[15], w08[15], w09[15], w10[15], w11[15], w12[15], w13[15], w14[15],
                                        S[14],   C[14]);
mips_wallace_unit wallace_unit15(s15, w00[15], w01[15], w02[15], w03[15], w04[15], w05[15], w06[15], w07[15], w08[15], w09[15], w10[15], w11[15], w12[15], w13[15], w14[15],
                                      w00[16], w01[16], w02[16], w03[16], w04[16], w05[16], w06[16], w07[16], w08[16], w09[16], w10[16], w11[16], w12[16], w13[16], w14[16],
                                        S[15],   C[15]);
mips_wallace_unit wallace_unit16(s16, w00[16], w01[16], w02[16], w03[16], w04[16], w05[16], w06[16], w07[16], w08[16], w09[16], w10[16], w11[16], w12[16], w13[16], w14[16],
                                      w00[17], w01[17], w02[17], w03[17], w04[17], w05[17], w06[17], w07[17], w08[17], w09[17], w10[17], w11[17], w12[17], w13[17], w14[17],
                                        S[16],   C[16]);
mips_wallace_unit wallace_unit17(s17, w00[17], w01[17], w02[17], w03[17], w04[17], w05[17], w06[17], w07[17], w08[17], w09[17], w10[17], w11[17], w12[17], w13[17], w14[17],
                                      w00[18], w01[18], w02[18], w03[18], w04[18], w05[18], w06[18], w07[18], w08[18], w09[18], w10[18], w11[18], w12[18], w13[18], w14[18],
                                        S[17],   C[17]);
mips_wallace_unit wallace_unit18(s18, w00[18], w01[18], w02[18], w03[18], w04[18], w05[18], w06[18], w07[18], w08[18], w09[18], w10[18], w11[18], w12[18], w13[18], w14[18],
                                      w00[19], w01[19], w02[19], w03[19], w04[19], w05[19], w06[19], w07[19], w08[19], w09[19], w10[19], w11[19], w12[19], w13[19], w14[19],
                                        S[18],   C[18]);
mips_wallace_unit wallace_unit19(s19, w00[19], w01[19], w02[19], w03[19], w04[19], w05[19], w06[19], w07[19], w08[19], w09[19], w10[19], w11[19], w12[19], w13[19], w14[19],
                                      w00[20], w01[20], w02[20], w03[20], w04[20], w05[20], w06[20], w07[20], w08[20], w09[20], w10[20], w11[20], w12[20], w13[20], w14[20],
                                        S[19],   C[19]);
mips_wallace_unit wallace_unit20(s20, w00[20], w01[20], w02[20], w03[20], w04[20], w05[20], w06[20], w07[20], w08[20], w09[20], w10[20], w11[20], w12[20], w13[20], w14[20],
                                      w00[21], w01[21], w02[21], w03[21], w04[21], w05[21], w06[21], w07[21], w08[21], w09[21], w10[21], w11[21], w12[21], w13[21], w14[21],
                                        S[20],   C[20]);
mips_wallace_unit wallace_unit21(s21, w00[21], w01[21], w02[21], w03[21], w04[21], w05[21], w06[21], w07[21], w08[21], w09[21], w10[21], w11[21], w12[21], w13[21], w14[21],
                                      w00[22], w01[22], w02[22], w03[22], w04[22], w05[22], w06[22], w07[22], w08[22], w09[22], w10[22], w11[22], w12[22], w13[22], w14[22],
                                        S[21],   C[21]);
mips_wallace_unit wallace_unit22(s22, w00[22], w01[22], w02[22], w03[22], w04[22], w05[22], w06[22], w07[22], w08[22], w09[22], w10[22], w11[22], w12[22], w13[22], w14[22],
                                      w00[23], w01[23], w02[23], w03[23], w04[23], w05[23], w06[23], w07[23], w08[23], w09[23], w10[23], w11[23], w12[23], w13[23], w14[23],
                                        S[22],   C[22]);
mips_wallace_unit wallace_unit23(s23, w00[23], w01[23], w02[23], w03[23], w04[23], w05[23], w06[23], w07[23], w08[23], w09[23], w10[23], w11[23], w12[23], w13[23], w14[23],
                                      w00[24], w01[24], w02[24], w03[24], w04[24], w05[24], w06[24], w07[24], w08[24], w09[24], w10[24], w11[24], w12[24], w13[24], w14[24],
                                        S[23],   C[23]);
mips_wallace_unit wallace_unit24(s24, w00[24], w01[24], w02[24], w03[24], w04[24], w05[24], w06[24], w07[24], w08[24], w09[24], w10[24], w11[24], w12[24], w13[24], w14[24],
                                      w00[25], w01[25], w02[25], w03[25], w04[25], w05[25], w06[25], w07[25], w08[25], w09[25], w10[25], w11[25], w12[25], w13[25], w14[25],
                                        S[24],   C[24]);
mips_wallace_unit wallace_unit25(s25, w00[25], w01[25], w02[25], w03[25], w04[25], w05[25], w06[25], w07[25], w08[25], w09[25], w10[25], w11[25], w12[25], w13[25], w14[25],
                                      w00[26], w01[26], w02[26], w03[26], w04[26], w05[26], w06[26], w07[26], w08[26], w09[26], w10[26], w11[26], w12[26], w13[26], w14[26],
                                        S[25],   C[25]);
mips_wallace_unit wallace_unit26(s26, w00[26], w01[26], w02[26], w03[26], w04[26], w05[26], w06[26], w07[26], w08[26], w09[26], w10[26], w11[26], w12[26], w13[26], w14[26],
                                      w00[27], w01[27], w02[27], w03[27], w04[27], w05[27], w06[27], w07[27], w08[27], w09[27], w10[27], w11[27], w12[27], w13[27], w14[27],
                                        S[26],   C[26]);
mips_wallace_unit wallace_unit27(s27, w00[27], w01[27], w02[27], w03[27], w04[27], w05[27], w06[27], w07[27], w08[27], w09[27], w10[27], w11[27], w12[27], w13[27], w14[27],
                                      w00[28], w01[28], w02[28], w03[28], w04[28], w05[28], w06[28], w07[28], w08[28], w09[28], w10[28], w11[28], w12[28], w13[28], w14[28],
                                        S[27],   C[27]);
mips_wallace_unit wallace_unit28(s28, w00[28], w01[28], w02[28], w03[28], w04[28], w05[28], w06[28], w07[28], w08[28], w09[28], w10[28], w11[28], w12[28], w13[28], w14[28],
                                      w00[29], w01[29], w02[29], w03[29], w04[29], w05[29], w06[29], w07[29], w08[29], w09[29], w10[29], w11[29], w12[29], w13[29], w14[29],
                                        S[28],   C[28]);
mips_wallace_unit wallace_unit29(s29, w00[29], w01[29], w02[29], w03[29], w04[29], w05[29], w06[29], w07[29], w08[29], w09[29], w10[29], w11[29], w12[29], w13[29], w14[29],
                                      w00[30], w01[30], w02[30], w03[30], w04[30], w05[30], w06[30], w07[30], w08[30], w09[30], w10[30], w11[30], w12[30], w13[30], w14[30],
                                        S[29],   C[29]);
mips_wallace_unit wallace_unit30(s30, w00[30], w01[30], w02[30], w03[30], w04[30], w05[30], w06[30], w07[30], w08[30], w09[30], w10[30], w11[30], w12[30], w13[30], w14[30],
                                      w00[31], w01[31], w02[31], w03[31], w04[31], w05[31], w06[31], w07[31], w08[31], w09[31], w10[31], w11[31], w12[31], w13[31], w14[31],
                                        S[30],   C[30]);
mips_wallace_unit wallace_unit31(s31, w00[31], w01[31], w02[31], w03[31], w04[31], w05[31], w06[31], w07[31], w08[31], w09[31], w10[31], w11[31], w12[31], w13[31], w14[31],
                                      w00[32], w01[32], w02[32], w03[32], w04[32], w05[32], w06[32], w07[32], w08[32], w09[32], w10[32], w11[32], w12[32], w13[32], w14[32],
                                        S[31],   C[31]);
mips_wallace_unit wallace_unit32(s32, w00[32], w01[32], w02[32], w03[32], w04[32], w05[32], w06[32], w07[32], w08[32], w09[32], w10[32], w11[32], w12[32], w13[32], w14[32],
                                      w00[33], w01[33], w02[33], w03[33], w04[33], w05[33], w06[33], w07[33], w08[33], w09[33], w10[33], w11[33], w12[33], w13[33], w14[33],
                                        S[32],   C[32]);
mips_wallace_unit wallace_unit33(s33, w00[33], w01[33], w02[33], w03[33], w04[33], w05[33], w06[33], w07[33], w08[33], w09[33], w10[33], w11[33], w12[33], w13[33], w14[33],
                                      w00[34], w01[34], w02[34], w03[34], w04[34], w05[34], w06[34], w07[34], w08[34], w09[34], w10[34], w11[34], w12[34], w13[34], w14[34],
                                        S[33],   C[33]);
mips_wallace_unit wallace_unit34(s34, w00[34], w01[34], w02[34], w03[34], w04[34], w05[34], w06[34], w07[34], w08[34], w09[34], w10[34], w11[34], w12[34], w13[34], w14[34],
                                      w00[35], w01[35], w02[35], w03[35], w04[35], w05[35], w06[35], w07[35], w08[35], w09[35], w10[35], w11[35], w12[35], w13[35], w14[35],
                                        S[34],   C[34]);
mips_wallace_unit wallace_unit35(s35, w00[35], w01[35], w02[35], w03[35], w04[35], w05[35], w06[35], w07[35], w08[35], w09[35], w10[35], w11[35], w12[35], w13[35], w14[35],
                                      w00[36], w01[36], w02[36], w03[36], w04[36], w05[36], w06[36], w07[36], w08[36], w09[36], w10[36], w11[36], w12[36], w13[36], w14[36],
                                        S[35],   C[35]);
mips_wallace_unit wallace_unit36(s36, w00[36], w01[36], w02[36], w03[36], w04[36], w05[36], w06[36], w07[36], w08[36], w09[36], w10[36], w11[36], w12[36], w13[36], w14[36],
                                      w00[37], w01[37], w02[37], w03[37], w04[37], w05[37], w06[37], w07[37], w08[37], w09[37], w10[37], w11[37], w12[37], w13[37], w14[37],
                                        S[36],   C[36]);
mips_wallace_unit wallace_unit37(s37, w00[37], w01[37], w02[37], w03[37], w04[37], w05[37], w06[37], w07[37], w08[37], w09[37], w10[37], w11[37], w12[37], w13[37], w14[37],
                                      w00[38], w01[38], w02[38], w03[38], w04[38], w05[38], w06[38], w07[38], w08[38], w09[38], w10[38], w11[38], w12[38], w13[38], w14[38],
                                        S[37],   C[37]);
mips_wallace_unit wallace_unit38(s38, w00[38], w01[38], w02[38], w03[38], w04[38], w05[38], w06[38], w07[38], w08[38], w09[38], w10[38], w11[38], w12[38], w13[38], w14[38],
                                      w00[39], w01[39], w02[39], w03[39], w04[39], w05[39], w06[39], w07[39], w08[39], w09[39], w10[39], w11[39], w12[39], w13[39], w14[39],
                                        S[38],   C[38]);
mips_wallace_unit wallace_unit39(s39, w00[39], w01[39], w02[39], w03[39], w04[39], w05[39], w06[39], w07[39], w08[39], w09[39], w10[39], w11[39], w12[39], w13[39], w14[39],
                                      w00[40], w01[40], w02[40], w03[40], w04[40], w05[40], w06[40], w07[40], w08[40], w09[40], w10[40], w11[40], w12[40], w13[40], w14[40],
                                        S[39],   C[39]);
mips_wallace_unit wallace_unit40(s40, w00[40], w01[40], w02[40], w03[40], w04[40], w05[40], w06[40], w07[40], w08[40], w09[40], w10[40], w11[40], w12[40], w13[40], w14[40],
                                      w00[41], w01[41], w02[41], w03[41], w04[41], w05[41], w06[41], w07[41], w08[41], w09[41], w10[41], w11[41], w12[41], w13[41], w14[41],
                                        S[40],   C[40]);
mips_wallace_unit wallace_unit41(s41, w00[41], w01[41], w02[41], w03[41], w04[41], w05[41], w06[41], w07[41], w08[41], w09[41], w10[41], w11[41], w12[41], w13[41], w14[41],
                                      w00[42], w01[42], w02[42], w03[42], w04[42], w05[42], w06[42], w07[42], w08[42], w09[42], w10[42], w11[42], w12[42], w13[42], w14[42],
                                        S[41],   C[41]);
mips_wallace_unit wallace_unit42(s42, w00[42], w01[42], w02[42], w03[42], w04[42], w05[42], w06[42], w07[42], w08[42], w09[42], w10[42], w11[42], w12[42], w13[42], w14[42],
                                      w00[43], w01[43], w02[43], w03[43], w04[43], w05[43], w06[43], w07[43], w08[43], w09[43], w10[43], w11[43], w12[43], w13[43], w14[43],
                                        S[42],   C[42]);
mips_wallace_unit wallace_unit43(s43, w00[43], w01[43], w02[43], w03[43], w04[43], w05[43], w06[43], w07[43], w08[43], w09[43], w10[43], w11[43], w12[43], w13[43], w14[43],
                                      w00[44], w01[44], w02[44], w03[44], w04[44], w05[44], w06[44], w07[44], w08[44], w09[44], w10[44], w11[44], w12[44], w13[44], w14[44],
                                        S[43],   C[43]);
mips_wallace_unit wallace_unit44(s44, w00[44], w01[44], w02[44], w03[44], w04[44], w05[44], w06[44], w07[44], w08[44], w09[44], w10[44], w11[44], w12[44], w13[44], w14[44],
                                      w00[45], w01[45], w02[45], w03[45], w04[45], w05[45], w06[45], w07[45], w08[45], w09[45], w10[45], w11[45], w12[45], w13[45], w14[45],
                                        S[44],   C[44]);
mips_wallace_unit wallace_unit45(s45, w00[45], w01[45], w02[45], w03[45], w04[45], w05[45], w06[45], w07[45], w08[45], w09[45], w10[45], w11[45], w12[45], w13[45], w14[45],
                                      w00[46], w01[46], w02[46], w03[46], w04[46], w05[46], w06[46], w07[46], w08[46], w09[46], w10[46], w11[46], w12[46], w13[46], w14[46],
                                        S[45],   C[45]);
mips_wallace_unit wallace_unit46(s46, w00[46], w01[46], w02[46], w03[46], w04[46], w05[46], w06[46], w07[46], w08[46], w09[46], w10[46], w11[46], w12[46], w13[46], w14[46],
                                      w00[47], w01[47], w02[47], w03[47], w04[47], w05[47], w06[47], w07[47], w08[47], w09[47], w10[47], w11[47], w12[47], w13[47], w14[47],
                                        S[46],   C[46]);
mips_wallace_unit wallace_unit47(s47, w00[47], w01[47], w02[47], w03[47], w04[47], w05[47], w06[47], w07[47], w08[47], w09[47], w10[47], w11[47], w12[47], w13[47], w14[47],
                                      w00[48], w01[48], w02[48], w03[48], w04[48], w05[48], w06[48], w07[48], w08[48], w09[48], w10[48], w11[48], w12[48], w13[48], w14[48],
                                        S[47],   C[47]);
mips_wallace_unit wallace_unit48(s48, w00[48], w01[48], w02[48], w03[48], w04[48], w05[48], w06[48], w07[48], w08[48], w09[48], w10[48], w11[48], w12[48], w13[48], w14[48],
                                      w00[49], w01[49], w02[49], w03[49], w04[49], w05[49], w06[49], w07[49], w08[49], w09[49], w10[49], w11[49], w12[49], w13[49], w14[49],
                                        S[48],   C[48]);
mips_wallace_unit wallace_unit49(s49, w00[49], w01[49], w02[49], w03[49], w04[49], w05[49], w06[49], w07[49], w08[49], w09[49], w10[49], w11[49], w12[49], w13[49], w14[49],
                                      w00[50], w01[50], w02[50], w03[50], w04[50], w05[50], w06[50], w07[50], w08[50], w09[50], w10[50], w11[50], w12[50], w13[50], w14[50],
                                        S[49],   C[49]);
mips_wallace_unit wallace_unit50(s50, w00[50], w01[50], w02[50], w03[50], w04[50], w05[50], w06[50], w07[50], w08[50], w09[50], w10[50], w11[50], w12[50], w13[50], w14[50],
                                      w00[51], w01[51], w02[51], w03[51], w04[51], w05[51], w06[51], w07[51], w08[51], w09[51], w10[51], w11[51], w12[51], w13[51], w14[51],
                                        S[50],   C[50]);
mips_wallace_unit wallace_unit51(s51, w00[51], w01[51], w02[51], w03[51], w04[51], w05[51], w06[51], w07[51], w08[51], w09[51], w10[51], w11[51], w12[51], w13[51], w14[51],
                                      w00[52], w01[52], w02[52], w03[52], w04[52], w05[52], w06[52], w07[52], w08[52], w09[52], w10[52], w11[52], w12[52], w13[52], w14[52],
                                        S[51],   C[51]);
mips_wallace_unit wallace_unit52(s52, w00[52], w01[52], w02[52], w03[52], w04[52], w05[52], w06[52], w07[52], w08[52], w09[52], w10[52], w11[52], w12[52], w13[52], w14[52],
                                      w00[53], w01[53], w02[53], w03[53], w04[53], w05[53], w06[53], w07[53], w08[53], w09[53], w10[53], w11[53], w12[53], w13[53], w14[53],
                                        S[52],   C[52]);
mips_wallace_unit wallace_unit53(s53, w00[53], w01[53], w02[53], w03[53], w04[53], w05[53], w06[53], w07[53], w08[53], w09[53], w10[53], w11[53], w12[53], w13[53], w14[53],
                                      w00[54], w01[54], w02[54], w03[54], w04[54], w05[54], w06[54], w07[54], w08[54], w09[54], w10[54], w11[54], w12[54], w13[54], w14[54],
                                        S[53],   C[53]);
mips_wallace_unit wallace_unit54(s54, w00[54], w01[54], w02[54], w03[54], w04[54], w05[54], w06[54], w07[54], w08[54], w09[54], w10[54], w11[54], w12[54], w13[54], w14[54],
                                      w00[55], w01[55], w02[55], w03[55], w04[55], w05[55], w06[55], w07[55], w08[55], w09[55], w10[55], w11[55], w12[55], w13[55], w14[55],
                                        S[54],   C[54]);
mips_wallace_unit wallace_unit55(s55, w00[55], w01[55], w02[55], w03[55], w04[55], w05[55], w06[55], w07[55], w08[55], w09[55], w10[55], w11[55], w12[55], w13[55], w14[55],
                                      w00[56], w01[56], w02[56], w03[56], w04[56], w05[56], w06[56], w07[56], w08[56], w09[56], w10[56], w11[56], w12[56], w13[56], w14[56],
                                        S[55],   C[55]);
mips_wallace_unit wallace_unit56(s56, w00[56], w01[56], w02[56], w03[56], w04[56], w05[56], w06[56], w07[56], w08[56], w09[56], w10[56], w11[56], w12[56], w13[56], w14[56],
                                      w00[57], w01[57], w02[57], w03[57], w04[57], w05[57], w06[57], w07[57], w08[57], w09[57], w10[57], w11[57], w12[57], w13[57], w14[57],
                                        S[56],   C[56]);
mips_wallace_unit wallace_unit57(s57, w00[57], w01[57], w02[57], w03[57], w04[57], w05[57], w06[57], w07[57], w08[57], w09[57], w10[57], w11[57], w12[57], w13[57], w14[57],
                                      w00[58], w01[58], w02[58], w03[58], w04[58], w05[58], w06[58], w07[58], w08[58], w09[58], w10[58], w11[58], w12[58], w13[58], w14[58],
                                        S[57],   C[57]);
mips_wallace_unit wallace_unit58(s58, w00[58], w01[58], w02[58], w03[58], w04[58], w05[58], w06[58], w07[58], w08[58], w09[58], w10[58], w11[58], w12[58], w13[58], w14[58],
                                      w00[59], w01[59], w02[59], w03[59], w04[59], w05[59], w06[59], w07[59], w08[59], w09[59], w10[59], w11[59], w12[59], w13[59], w14[59],
                                        S[58],   C[58]);
mips_wallace_unit wallace_unit59(s59, w00[59], w01[59], w02[59], w03[59], w04[59], w05[59], w06[59], w07[59], w08[59], w09[59], w10[59], w11[59], w12[59], w13[59], w14[59],
                                      w00[60], w01[60], w02[60], w03[60], w04[60], w05[60], w06[60], w07[60], w08[60], w09[60], w10[60], w11[60], w12[60], w13[60], w14[60],
                                        S[59],   C[59]);
mips_wallace_unit wallace_unit60(s60, w00[60], w01[60], w02[60], w03[60], w04[60], w05[60], w06[60], w07[60], w08[60], w09[60], w10[60], w11[60], w12[60], w13[60], w14[60],
                                      w00[61], w01[61], w02[61], w03[61], w04[61], w05[61], w06[61], w07[61], w08[61], w09[61], w10[61], w11[61], w12[61], w13[61], w14[61],
                                        S[60],   C[60]);
mips_wallace_unit wallace_unit61(s61, w00[61], w01[61], w02[61], w03[61], w04[61], w05[61], w06[61], w07[61], w08[61], w09[61], w10[61], w11[61], w12[61], w13[61], w14[61],
                                      w00[62], w01[62], w02[62], w03[62], w04[62], w05[62], w06[62], w07[62], w08[62], w09[62], w10[62], w11[62], w12[62], w13[62], w14[62],
                                        S[61],   C[61]);
mips_wallace_unit wallace_unit62(s62, w00[62], w01[62], w02[62], w03[62], w04[62], w05[62], w06[62], w07[62], w08[62], w09[62], w10[62], w11[62], w12[62], w13[62], w14[62],
                                      w00[63], w01[63], w02[63], w03[63], w04[63], w05[63], w06[63], w07[63], w08[63], w09[63], w10[63], w11[63], w12[63], w13[63], w14[63],
                                        S[62],   C[62]);
mips_wallace_unit wallace_unit63(s63, w00[63], w01[63], w02[63], w03[63], w04[63], w05[63], w06[63], w07[63], w08[63], w09[63], w10[63], w11[63], w12[63], w13[63], w14[63],
                                      w00[64], w01[64], w02[64], w03[64], w04[64], w05[64], w06[64], w07[64], w08[64], w09[64], w10[64], w11[64], w12[64], w13[64], w14[64],
                                        S[63],   C[63]);
mips_wallace_unit wallace_unit64(s64, w00[64], w01[64], w02[64], w03[64], w04[64], w05[64], w06[64], w07[64], w08[64], w09[64], w10[64], w11[64], w12[64], w13[64], w14[64],
                                      w00[65], w01[65], w02[65], w03[65], w04[65], w05[65], w06[65], w07[65], w08[65], w09[65], w10[65], w11[65], w12[65], w13[65], w14[65],
                                        S[64],   C[64]);
mips_wallace_unit wallace_unit65(s65, w00[65], w01[65], w02[65], w03[65], w04[65], w05[65], w06[65], w07[65], w08[65], w09[65], w10[65], w11[65], w12[65], w13[65], w14[65],
                                      w00[66], w01[66], w02[66], w03[66], w04[66], w05[66], w06[66], w07[66], w08[66], w09[66], w10[66], w11[66], w12[66], w13[66], w14[66],
                                        S[65],   C[65]);

mips_booth_stage booth_stage(A, B, p00, p01, p02, p03, p04, p05, p06, p07, p08, p09, p10, p11, p12, p13, p14, p15, p16,
                                   C00, C01, C02, C03, C04, C05, C06, C07, C08, C09, C10, C11, C12, C13, C14, C15, C16);
endmodule


module mips_booth_stage (
    input  wire [32:0] A,
    input  wire [32:0] B,
    output wire [65:0] p00, p01, p02, p03, p04, p05, 
    output wire [65:0] p06, p07, p08, p09, p10, p11,
    output wire [65:0] p12, p13, p14, p15, p16,
    output wire        C00, C01, C02, C03, C04, C05, 
    output wire        C06, C07, C08, C09, C10, C11, 
    output wire        C12, C13, C14, C15, C16
    );

wire [34:0] booth_B  = {B[32], B, 1'b0};
wire [65:0] booth_p00, booth_p01, booth_p02, booth_p03, booth_p04, booth_p05, booth_p06, booth_p07, booth_p08, booth_p09;
wire [65:0] booth_p10, booth_p11, booth_p12, booth_p13, booth_p14, booth_p15, booth_p16;

assign p00 = {booth_p00[65:0]       };
assign p01 = {booth_p01[63:0],  2'd0};
assign p02 = {booth_p02[61:0],  4'd0};
assign p03 = {booth_p03[59:0],  6'd0};
assign p04 = {booth_p04[57:0],  8'd0};
assign p05 = {booth_p05[55:0], 10'd0};
assign p06 = {booth_p06[53:0], 12'd0};
assign p07 = {booth_p07[51:0], 14'd0};
assign p08 = {booth_p08[49:0], 16'd0};
assign p09 = {booth_p09[47:0], 18'd0};
assign p10 = {booth_p10[45:0], 20'd0};
assign p11 = {booth_p11[43:0], 22'd0};
assign p12 = {booth_p12[41:0], 24'd0};
assign p13 = {booth_p13[39:0], 26'd0};
assign p14 = {booth_p14[37:0], 28'd0};
assign p15 = {booth_p15[35:0], 30'd0};
assign p16 = {booth_p16[33:0], 32'd0};

mips_booth_unit both_unit00(A, booth_B[ 2: 0], booth_p00, C00);
mips_booth_unit both_unit01(A, booth_B[ 4: 2], booth_p01, C01);
mips_booth_unit both_unit02(A, booth_B[ 6: 4], booth_p02, C02);
mips_booth_unit both_unit03(A, booth_B[ 8: 6], booth_p03, C03);
mips_booth_unit both_unit04(A, booth_B[10: 8], booth_p04, C04);
mips_booth_unit both_unit05(A, booth_B[12:10], booth_p05, C05);
mips_booth_unit both_unit06(A, booth_B[14:12], booth_p06, C06);
mips_booth_unit both_unit07(A, booth_B[16:14], booth_p07, C07);
mips_booth_unit both_unit08(A, booth_B[18:16], booth_p08, C08);
mips_booth_unit both_unit09(A, booth_B[20:18], booth_p09, C09);
mips_booth_unit both_unit10(A, booth_B[22:20], booth_p10, C10);
mips_booth_unit both_unit11(A, booth_B[24:22], booth_p11, C11);
mips_booth_unit both_unit12(A, booth_B[26:24], booth_p12, C12);
mips_booth_unit both_unit13(A, booth_B[28:26], booth_p13, C13);
mips_booth_unit both_unit14(A, booth_B[30:28], booth_p14, C14);
mips_booth_unit both_unit15(A, booth_B[32:30], booth_p15, C15);
mips_booth_unit both_unit16(A, booth_B[34:32], booth_p16, C16);

endmodule

module mips_booth_unit (
    input  wire [32:0] A,
    input  wire [ 2:0] B,
    output wire [65:0] P,
    output wire        C
    );

wire [32:0] Ac = (~A) + 33'd1;

assign {P, C} = ({67{B == 3'b001}} & {{33{A [32]}}, A , 1'b0 })
              | ({67{B == 3'b010}} & {{33{A [32]}}, A , 1'b0 })
              | ({67{B == 3'b011}} & {{32{A [32]}}, A , 2'b00})
              | ({67{B == 3'b100}} & {{32{Ac[32]}}, Ac, 2'b00})
              | ({67{B == 3'b101}} & {{33{Ac[32]}}, Ac, 1'b0 })
              | ({67{B == 3'b110}} & {{33{Ac[32]}}, Ac, 1'b0 });

endmodule


module mips_add_carry (
    input  wire A,
    input  wire B,
    input  wire D,
    output wire S,
    output wire C
    );

assign S = A ^ B ^ D;
assign C = (A & B) | (A & D) | (B & D);

endmodule


module mips_wallace_unit (
    input  wire [16:0] s,
    input  wire        in_00 , in_01 , in_02 , in_03 , in_04 ,
    input  wire        in_05 , in_06 , in_07 , in_08 , in_09 ,
    input  wire        in_10 , in_11 , in_12 , in_13 , in_14 ,
    output wire        out_00, out_01, out_02, out_03, out_04,
    output wire        out_05, out_06, out_07, out_08, out_09,
    output wire        out_10, out_11, out_12, out_13, out_14,
    output wire        S,
    output wire        C
);

wire w00, w01, w02, w03, w04, w05, w06, w07, w08, w09, w10, w11, w12, w13, w14;

mips_add_carry add_carry00( s[ 1],  s[ 0],  1'b0 , w00, out_00);
mips_add_carry add_carry01( s[ 4],  s[ 3],  s[ 2], w01, out_01);
mips_add_carry add_carry02( s[ 7],  s[ 6],  s[ 5], w02, out_02);
mips_add_carry add_carry03( s[10],  s[ 9],  s[ 8], w03, out_03);
mips_add_carry add_carry04( s[13],  s[12],  s[11], w04, out_04);
mips_add_carry add_carry05( s[16],  s[15],  s[14], w05, out_05);

mips_add_carry add_carry06( in_02,  in_01,  in_00, w06, out_06);
mips_add_carry add_carry07( in_05,  in_04,  in_03, w07, out_07);
mips_add_carry add_carry08(   w02,    w01,    w00, w08, out_08);
mips_add_carry add_carry09(   w05,    w04,    w03, w09, out_09);

mips_add_carry add_carry10(   w06,  in_07,  in_06, w10, out_10);
mips_add_carry add_carry11(   w09,    w08,    w07, w11, out_11);

mips_add_carry add_carry12( in_10,  in_09,  in_08, w12, out_12);
mips_add_carry add_carry13(   w11,    w10,  in_11, w13, out_13);

mips_add_carry add_carry14(   w13,    w12,  in_12, w14, out_14);

mips_add_carry add_carry15(   w14,  in_14,  in_13,   S,      C);

endmodule
